module tt_um_and(
  input logic clk,
  input logic reset,
  input logic [7:0] a, b,
  output logic [7:0] Y
);
  
  assign Y = a & b;
endmodule
